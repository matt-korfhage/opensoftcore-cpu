library ieee; use ieee.std_logic_1164.all; 
package dseg7font is  
 
  constant dseg7_0:    std_logic_vector(7 downto 0) := B"11000000";  
  constant dseg7_1:    std_logic_vector(7 downto 0) := B"11111001";  
  constant dseg7_2:    std_logic_vector(7 downto 0) := B"10100100";  
  constant dseg7_3:    std_logic_vector(7 downto 0) := B"10110000";  
  constant dseg7_4:    std_logic_vector(7 downto 0) := B"10011001"; --Completed 
  constant dseg7_5:    std_logic_vector(7 downto 0) := B"10010010"; 
  constant dseg7_6:    std_logic_vector(7 downto 0) := B"10000010"; 
  constant dseg7_7:    std_logic_vector(7 downto 0) := B"11011000"; 
  constant dseg7_8:    std_logic_vector(7 downto 0) := B"10000000"; 
  constant dseg7_9:    std_logic_vector(7 downto 0) := B"10010000"; 
  constant dseg7_a:    std_logic_vector(7 downto 0) := B"10001000"; 
  constant dseg7_b:    std_logic_vector(7 downto 0) := B"10000011"; 
  constant dseg7_c:    std_logic_vector(7 downto 0) := B"10100111"; 
  constant dseg7_d:    std_logic_vector(7 downto 0) := B"10100001"; --Completed 
  constant dseg7_e:    std_logic_vector(7 downto 0) := B"10000110"; --Completed  
  constant dseg7_f:    std_logic_vector(7 downto 0) := B"10001110"; 
  constant dseg7_g:    std_logic_vector(7 downto 0) := B"11000010"; --Completed
  constant dseg7_h:    std_logic_vector(7 downto 0) := B"10001011"; 
  constant dseg7_i:    std_logic_vector(7 downto 0) := B"11111011"; 
  constant dseg7_j:    std_logic_vector(7 downto 0) := B"11100001"; 
  constant dseg7_k:    std_logic_vector(7 downto 0) := B"10001010"; 
  constant dseg7_l:    std_logic_vector(7 downto 0) := B"11000111"; 
  constant dseg7_m:    std_logic_vector(7 downto 0) := B"11001000";  
  constant dseg7_n:    std_logic_vector(7 downto 0) := B"10101011"; --Completed 
  constant dseg7_o:    std_logic_vector(7 downto 0) := B"10100011"; 
  constant dseg7_p:    std_logic_vector(7 downto 0) := B"10001100"; 
  constant dseg7_q:    std_logic_vector(7 downto 0) := B"10011000"; 
  constant dseg7_r:    std_logic_vector(7 downto 0) := B"10101111"; --Completed
  constant dseg7_s:    std_logic_vector(7 downto 0) := B"10010010"; 
  constant dseg7_t:    std_logic_vector(7 downto 0) := B"10000111"; 
  constant dseg7_u:    std_logic_vector(7 downto 0) := B"11100011"; --Completed 
  constant dseg7_v:    std_logic_vector(7 downto 0) := B"11000001"; 
  constant dseg7_w:    std_logic_vector(7 downto 0) := B"10000001"; --Completed 
  constant dseg7_x:    std_logic_vector(7 downto 0) := B"10001001"; --Completed
  constant dseg7_y:    std_logic_vector(7 downto 0) := B"10010001"; 
  constant dseg7_z:    std_logic_vector(7 downto 0) := B"11100100"; 
  constant dseg7_blank:std_logic_vector(7 downto 0) := B"11111111"; 
  
  end package dseg7font;	